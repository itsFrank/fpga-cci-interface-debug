// SCFIFO.v 

// Generated using ACDS version 16.0 211
`timescale 1 ps / 1 ps
module SCFIFO #(
	parameter FWFT = "OFF",
	parameter DATA_WIDTH = 512,
	parameter DEPTH = 64,
	parameter COUNT_WIDTH = 6,
	parameter ALM_FULL_DIFF = 0,
	parameter ALM_EMPTY_DIFF = 0
)
(
	input  wire         clock, 
	i_fifo.to_fifo 		fifo_if
);

	localparam ALM_FULL_VALUE = DEPTH - ALM_FULL_DIFF;

	scfifo  scfifo_component (
		.clock (clock),
		.data  (fifo_if.data_in),  
		.rdreq (fifo_if.rd_en), 
		.sclr  (fifo_if.reset),  
		.wrreq (fifo_if.wr_en), 
		.empty (fifo_if.empty),  
		.full  (fifo_if.full),  
		.q     (fifo_if.data_out),     
		.usedw (fifo_if.count),
		.aclr (),
		.almost_empty (fifo_if.alm_empty),
		.almost_full (fifo_if.alm_full),
		.eccstatus ()
	);
	defparam
		scfifo_component.add_ram_output_register  = "ON",
		scfifo_component.enable_ecc  = "FALSE",
		scfifo_component.intended_device_family  = "Arria 10",
		scfifo_component.lpm_numwords  = DEPTH,
		scfifo_component.lpm_showahead  = FWFT,
		scfifo_component.lpm_type  = "scfifo",
		scfifo_component.lpm_width  = DATA_WIDTH,
		scfifo_component.lpm_widthu  = COUNT_WIDTH,
		scfifo_component.overflow_checking  = "OFF",
		scfifo_component.underflow_checking  = "OFF",
		scfifo_component.almost_empty_value  = ALM_EMPTY_DIFF, 
		scfifo_component.almost_full_value  = ALM_FULL_VALUE,
		scfifo_component.use_eab  = "ON";
endmodule